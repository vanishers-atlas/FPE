library ieee;
use ieee.std_logic_1164.all;

entity testbench is

end entity;

architecture arch of testbench is
	signal 	clock : std_logic := '0';
	signal	kickoff : std_logic := '0';
	signal	running : std_logic;

	signal	PUT_FIFO_0_data  : std_logic_vector(39 downto 0);
	signal	PUT_FIFO_0_write : std_logic;
begin
  UUT : entity work.test_FPE_inst(arch)
		port map (
			PUT_FIFO_0_data  => PUT_FIFO_0_data,
			PUT_FIFO_0_write => PUT_FIFO_0_write,
			clock => clock,
			kickoff => kickoff,
			running => running
		);

	-- Clock generate process
	clock_gen : process
	begin
	  loop
	    clock <= not clock;
	    wait for 50 ns;
	  end loop;
	end process;

	-- Signal kickoff after 200 ns
	kickoff <= '1' after 200 ns, '0' after 300 ns;


	spoff_PUT_FIFO_0 : process
	  variable  data_index : integer := 0;
	  type  data_array is array (0 to 223) of std_logic_vector(39 downto 0);
	  constant test_data : data_array :=
	  (
			-- Test MOV and ACC persistances
			"0000000000000000000000000000000000000000", "0000000000000000000000000000000000000000",
			"0000000000000000000011111111111111111111", "0000000000000000000011111111111111111111",
			"1111111111111111111100000000000000000000", "1111111111111111111100000000000000000000",
			"1111111111111111111111111111111111111111", "1111111111111111111111111111111111111111",

			-- Test LSH 1
			"0010001000100010001000100010001000100010", "0100010001000100010001000100010001000100",
			"1000100010001000100010001000100010001000", "0001000100010001000100010001000100010000",
			"0100010001000100010001000100010001000100", "1000100010001000100010001000100010001000",
			"0001000100010001000100010001000100010000", "0010001000100010001000100010001000100000",
			"1000100010001000100010001000100010001000", "0001000100010001000100010001000100010000",
			"0010001000100010001000100010001000100000", "0100010001000100010001000100010001000000",
			"0001000100010001000100010001000100010000", "0010001000100010001000100010001000100000",
			"0100010001000100010001000100010001000000", "1000100010001000100010001000100010000000",

			-- Test LSH 2
			"0100010001000100010001000100010001000100", "0001000100010001000100010001000100010000",
			"0100010001000100010001000100010001000000", "0001000100010001000100010001000100000000",
			"1000100010001000100010001000100010001000", "0010001000100010001000100010001000100000",
			"1000100010001000100010001000100010000000", "0010001000100010001000100010001000000000",
			"0001000100010001000100010001000100010000", "0100010001000100010001000100010001000000",
			"0001000100010001000100010001000100000000", "0100010001000100010001000100010000000000",
			"0010001000100010001000100010001000100000", "1000100010001000100010001000100010000000",
			"0010001000100010001000100010001000000000", "1000100010001000100010001000100000000000",

			-- Test LSH 3
			"1000100010001000100010001000100010001000", "0100010001000100010001000100010001000000",
			"0010001000100010001000100010001000000000", "0001000100010001000100010001000000000000",
			"0001000100010001000100010001000100010000", "1000100010001000100010001000100010000000",
			"0100010001000100010001000100010000000000", "0010001000100010001000100010000000000000",
			"0010001000100010001000100010001000100000", "0001000100010001000100010001000100000000",
			"1000100010001000100010001000100000000000", "0100010001000100010001000100000000000000",
			"0100010001000100010001000100010001000000", "0010001000100010001000100010001000000000",
			"0001000100010001000100010001000000000000", "1000100010001000100010001000000000000000",

			-- Test LRL 1
			"0010001000100010001000100010001000100010", "0100010001000100010001000100010001000100",
			"1000100010001000100010001000100010001000", "0001000100010001000100010001000100010001",
			"0100010001000100010001000100010001000100", "1000100010001000100010001000100010001000",
			"0001000100010001000100010001000100010001", "0010001000100010001000100010001000100010",
			"1000100010001000100010001000100010001000", "0001000100010001000100010001000100010001",
			"0010001000100010001000100010001000100010", "0100010001000100010001000100010001000100",
			"0001000100010001000100010001000100010001", "0010001000100010001000100010001000100010",
			"0100010001000100010001000100010001000100", "1000100010001000100010001000100010001000",

			-- Test LRL 2
			"0100010001000100010001000100010001000100", "0001000100010001000100010001000100010001",
			"0100010001000100010001000100010001000100", "0001000100010001000100010001000100010001",
			"1000100010001000100010001000100010001000", "0010001000100010001000100010001000100010",
			"1000100010001000100010001000100010001000", "0010001000100010001000100010001000100010",
			"0001000100010001000100010001000100010001", "0100010001000100010001000100010001000100",
			"0001000100010001000100010001000100010001", "0100010001000100010001000100010001000100",
			"0010001000100010001000100010001000100010", "1000100010001000100010001000100010001000",
			"0010001000100010001000100010001000100010", "1000100010001000100010001000100010001000",

			-- Test LRL 3
			"1000100010001000100010001000100010001000", "0100010001000100010001000100010001000100",
			"0010001000100010001000100010001000100010", "0001000100010001000100010001000100010001",
			"0001000100010001000100010001000100010001", "1000100010001000100010001000100010001000",
			"0100010001000100010001000100010001000100", "0010001000100010001000100010001000100010",
			"0010001000100010001000100010001000100010", "0001000100010001000100010001000100010001",
			"1000100010001000100010001000100010001000", "0100010001000100010001000100010001000100",
			"0100010001000100010001000100010001000100", "0010001000100010001000100010001000100010",
			"0001000100010001000100010001000100010001", "1000100010001000100010001000100010001000",

			-- Test RSH 1
			"0100010001000100010001000100010001000100", "0010001000100010001000100010001000100010",
			"0001000100010001000100010001000100010001", "0000100010001000100010001000100010001000",
			"0010001000100010001000100010001000100010", "0001000100010001000100010001000100010001",
			"0000100010001000100010001000100010001000", "0000010001000100010001000100010001000100",
			"0001000100010001000100010001000100010001", "0000100010001000100010001000100010001000",
			"0000010001000100010001000100010001000100", "0000001000100010001000100010001000100010",
			"0000100010001000100010001000100010001000", "0000010001000100010001000100010001000100",
			"0000001000100010001000100010001000100010", "0000000100010001000100010001000100010001",

			-- Test RSH 2
			"0010001000100010001000100010001000100010", "0000100010001000100010001000100010001000",
			"0000001000100010001000100010001000100010", "0000000010001000100010001000100010001000",
			"0001000100010001000100010001000100010001", "0000010001000100010001000100010001000100",
			"0000000100010001000100010001000100010001", "0000000001000100010001000100010001000100",
			"0000100010001000100010001000100010001000", "0000001000100010001000100010001000100010",
			"0000000010001000100010001000100010001000", "0000000000100010001000100010001000100010",
			"0000010001000100010001000100010001000100", "0000000100010001000100010001000100010001",
			"0000000001000100010001000100010001000100", "0000000000010001000100010001000100010001",

			-- Test RSH 3
			"0001000100010001000100010001000100010001", "0000001000100010001000100010001000100010",
			"0000000001000100010001000100010001000100", "0000000000001000100010001000100010001000",

			"0000100010001000100010001000100010001000", "0000000100010001000100010001000100010001",
			"0000000000100010001000100010001000100010", "0000000000000100010001000100010001000100",

			"0000010001000100010001000100010001000100", "0000000010001000100010001000100010001000",
			"0000000000010001000100010001000100010001", "0000000000000010001000100010001000100010",

			"0000001000100010001000100010001000100010", "0000000001000100010001000100010001000100",
			"0000000000001000100010001000100010001000", "0000000000000001000100010001000100010001",

			-- Test RRL 1
			"0100010001000100010001000100010001000100", "0010001000100010001000100010001000100010",
			"0001000100010001000100010001000100010001", "1000100010001000100010001000100010001000",
			"0010001000100010001000100010001000100010", "0001000100010001000100010001000100010001",
			"1000100010001000100010001000100010001000", "0100010001000100010001000100010001000100",
			"0001000100010001000100010001000100010001", "1000100010001000100010001000100010001000",
			"0100010001000100010001000100010001000100", "0010001000100010001000100010001000100010",
			"1000100010001000100010001000100010001000", "0100010001000100010001000100010001000100",
			"0010001000100010001000100010001000100010", "0001000100010001000100010001000100010001",

			-- Test RRL 2
			"0010001000100010001000100010001000100010", "1000100010001000100010001000100010001000",
			"0010001000100010001000100010001000100010", "1000100010001000100010001000100010001000",
			"0001000100010001000100010001000100010001", "0100010001000100010001000100010001000100",
			"0001000100010001000100010001000100010001", "0100010001000100010001000100010001000100",
			"1000100010001000100010001000100010001000", "0010001000100010001000100010001000100010",
			"1000100010001000100010001000100010001000", "0010001000100010001000100010001000100010",
			"0100010001000100010001000100010001000100", "0001000100010001000100010001000100010001",
			"0100010001000100010001000100010001000100", "0001000100010001000100010001000100010001",

			-- Test RRL 3
			"0001000100010001000100010001000100010001", "0010001000100010001000100010001000100010",
			"0100010001000100010001000100010001000100", "1000100010001000100010001000100010001000",
			"1000100010001000100010001000100010001000", "0001000100010001000100010001000100010001",
			"0010001000100010001000100010001000100010", "0100010001000100010001000100010001000100",
			"0100010001000100010001000100010001000100", "1000100010001000100010001000100010001000",
			"0001000100010001000100010001000100010001", "0010001000100010001000100010001000100010",
			"0010001000100010001000100010001000100010", "0100010001000100010001000100010001000100",
			"1000100010001000100010001000100010001000", "0001000100010001000100010001000100010001",

			-- Test NOT
			"1111111111111111111111111111111111111111", "0000000000000000000000000000000000000000",
			"1111111111111111111100000000000000000000", "0000000000000000000011111111111111111111",
			"0000000000000000000011111111111111111111", "1111111111111111111100000000000000000000",
			"0000000000000000000000000000000000000000", "1111111111111111111111111111111111111111",

			-- Test MUL
			"0000000000000000000000000000000000000000", "0000000000000000000000000000000000000000",
			"0000000000000000000000000000000000000001", "0000000000000000000011111110111100000001",
			"0000000000000000000000000000000000000000", "0000000000000000000000000000000000000000",
			"0000000000000000000000000000000000000001", "0000000000000000000011111110111100000001",
			"0000000000000000000000000000000000000000", "0000000000000000000000000000000000000000",
			"0000000000000000000000000000000000000001", "0000000000000000000011111110111100000001",
			"0000000000000000000000000000000000000000", "0000000000000000000000000000000000000001",
			"0000000000000000000000000000000000000100", "0000000000000000000000001111111000000001"
	  );
	begin
	  wait until running = '1';

	  -- Happen expected output
	  while 0 <= data_index and data_index < test_data'Length loop

	    wait until rising_edge(clock) and PUT_FIFO_0_write = '1';

	    -- Check the data is correct
	    assert(PUT_FIFO_0_data = test_data(data_index))
	      report "PUT_FIFO_0: Incorrect " & integer'Image(data_index) & " th output"
	      severity error;
	    assert(PUT_FIFO_0_data /= test_data(data_index))
	      report "PUT_FIFO_0: Correct " & integer'Image(data_index) & " th output"
	      severity note;

	      -- Advance to output index
	      data_index := data_index + 1;
	  end loop;

	  -- Mark all expected output given
	  report "PUT_FIFO_0: All expected output received" severity note;

	  -- Check for unexpected output
	  loop
	    wait until rising_edge(clock) and PUT_FIFO_0_write = '1';
	    report "PUT_FIFO_0: Extra output" severity error;
	  end loop;

	end process;

end architecture;
