library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

package ssp_instencoding is
  constant NOP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(0, 4));
  constant ADDMULSRA_MMIM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(1, 4));
  constant ADDMULSRA_MPIP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(2, 4));
  constant ADDMULSRA_FMIM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(3, 4));
  constant SUBMULSRA_MMIM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(4, 4));
  constant SUBMULSRA_MFIF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(5, 4));
  constant SUBMULSRA_FMIM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(6, 4));
  constant JMP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(7, 4));
  constant SETSMRB_0 : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(8, 4));
  constant ADDMUL_RRRR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMUL_RRRM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMUL_RRRI : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMUL_RRRF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMUL_RRRP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMUL_RRMR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMUL_RRMM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMUL_RRMI : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMUL_RRMF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMUL_RRMP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMUL_RRIR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMUL_RRIM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMUL_RRIF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMUL_RRIP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMUL_RRFR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMUL_RRFM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMUL_RRFI : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMUL_RRFF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMUL_RRFP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMUL_RRPR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMUL_RRPM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMUL_RRPI : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMUL_RRPF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMUL_RRPP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMUL_RMRR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMUL_RMRM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMUL_RMRI : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMUL_RMRF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMUL_RMRP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMUL_RMMR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMUL_RMMI : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMUL_RMMF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMUL_RMMP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMUL_RMIR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMUL_RMIM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMUL_RMIF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMUL_RMIP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMUL_RMFR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMUL_RMFM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMUL_RMFI : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMUL_RMFF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMUL_RMFP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMUL_RMPR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMUL_RMPM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMUL_RMPI : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMUL_RMPF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMUL_RMPP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMUL_RIRR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMUL_RIRM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMUL_RIRF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMUL_RIRP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMUL_RIMR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMUL_RIMM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMUL_RIMF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMUL_RIMP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMUL_RIFR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMUL_RIFM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMUL_RIFF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMUL_RIFP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMUL_RIPR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMUL_RIPM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMUL_RIPF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMUL_RIPP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMUL_RFRR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMUL_RFRM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMUL_RFRI : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMUL_RFRF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMUL_RFRP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMUL_RFMR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMUL_RFMM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMUL_RFMI : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMUL_RFMF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMUL_RFMP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMUL_RFIR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMUL_RFIM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMUL_RFIF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMUL_RFIP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMUL_RFFR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMUL_RFFM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMUL_RFFI : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMUL_RFPR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMUL_RFPM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMUL_RFPI : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMUL_RPRR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMUL_RPRM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMUL_RPRI : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMUL_RPRF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMUL_RPRP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMUL_RPMR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMUL_RPMM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMUL_RPMI : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMUL_RPMF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMUL_RPMP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMUL_RPIR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMUL_RPIM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMUL_RPIF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMUL_RPIP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMUL_RPFR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMUL_RPFM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMUL_RPFI : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMUL_RPPR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMUL_RPPM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMUL_RPPI : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMUL_MRRR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMUL_MRRM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMUL_MRRI : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMUL_MRRF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMUL_MRRP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMUL_MRMR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMUL_MRMM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMUL_MRMI : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMUL_MRMF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMUL_MRMP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMUL_MRIR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMUL_MRIM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMUL_MRIF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMUL_MRIP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMUL_MRFR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMUL_MRFM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMUL_MRFI : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMUL_MRFF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMUL_MRFP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMUL_MRPR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMUL_MRPM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMUL_MRPI : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMUL_MRPF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMUL_MRPP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMUL_MMRR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMUL_MMRM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMUL_MMRI : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMUL_MMRF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMUL_MMRP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMUL_MMMR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMUL_MMMI : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMUL_MMMF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMUL_MMMP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMUL_MMIR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMUL_MMIM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMUL_MMIF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMUL_MMIP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMUL_MMFR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMUL_MMFM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMUL_MMFI : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMUL_MMFF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMUL_MMFP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMUL_MMPR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMUL_MMPM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMUL_MMPI : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMUL_MMPF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMUL_MMPP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMUL_MIRR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMUL_MIRM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMUL_MIRF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMUL_MIRP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMUL_MIMR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMUL_MIMM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMUL_MIMF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMUL_MIMP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMUL_MIFR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMUL_MIFM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMUL_MIFF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMUL_MIFP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMUL_MIPR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMUL_MIPM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMUL_MIPF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMUL_MIPP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMUL_MFRR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMUL_MFRM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMUL_MFRI : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMUL_MFRF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMUL_MFRP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMUL_MFMR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMUL_MFMM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMUL_MFMI : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMUL_MFMF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMUL_MFMP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMUL_MFIR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMUL_MFIM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMUL_MFIF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMUL_MFIP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMUL_MFFR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMUL_MFFM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMUL_MFFI : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMUL_MFPR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMUL_MFPM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMUL_MFPI : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMUL_MPRR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMUL_MPRM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMUL_MPRI : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMUL_MPRF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMUL_MPRP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMUL_MPMR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMUL_MPMM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMUL_MPMI : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMUL_MPMF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMUL_MPMP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMUL_MPIR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMUL_MPIM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMUL_MPIF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMUL_MPIP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMUL_MPFR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMUL_MPFM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMUL_MPFI : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMUL_MPPR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMUL_MPPM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMUL_MPPI : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMUL_FRRR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMUL_FRRM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMUL_FRRI : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMUL_FRRF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMUL_FRRP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMUL_FRMR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMUL_FRMM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMUL_FRMI : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMUL_FRMF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMUL_FRMP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMUL_FRIR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMUL_FRIM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMUL_FRIF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMUL_FRIP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMUL_FRFR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMUL_FRFM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMUL_FRFI : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMUL_FRFF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMUL_FRFP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMUL_FRPR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMUL_FRPM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMUL_FRPI : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMUL_FRPF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMUL_FRPP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMUL_FMRR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMUL_FMRM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMUL_FMRI : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMUL_FMRF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMUL_FMRP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMUL_FMMR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMUL_FMMI : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMUL_FMMF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMUL_FMMP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMUL_FMIR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMUL_FMIM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMUL_FMIF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMUL_FMIP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMUL_FMFR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMUL_FMFM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMUL_FMFI : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMUL_FMFF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMUL_FMFP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMUL_FMPR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMUL_FMPM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMUL_FMPI : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMUL_FMPF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMUL_FMPP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMUL_FIRR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMUL_FIRM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMUL_FIRF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMUL_FIRP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMUL_FIMR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMUL_FIMM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMUL_FIMF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMUL_FIMP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMUL_FIFR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMUL_FIFM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMUL_FIFF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMUL_FIFP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMUL_FIPR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMUL_FIPM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMUL_FIPF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMUL_FIPP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMUL_FFRR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMUL_FFRM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMUL_FFRI : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMUL_FFRF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMUL_FFRP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMUL_FFMR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMUL_FFMM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMUL_FFMI : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMUL_FFMF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMUL_FFMP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMUL_FFIR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMUL_FFIM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMUL_FFIF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMUL_FFIP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMUL_FFFR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMUL_FFFM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMUL_FFFI : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMUL_FFPR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMUL_FFPM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMUL_FFPI : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMUL_FPRR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMUL_FPRM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMUL_FPRI : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMUL_FPRF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMUL_FPRP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMUL_FPMR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMUL_FPMM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMUL_FPMI : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMUL_FPMF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMUL_FPMP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMUL_FPIR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMUL_FPIM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMUL_FPIF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMUL_FPIP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMUL_FPFR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMUL_FPFM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMUL_FPFI : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMUL_FPPR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMUL_FPPM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMUL_FPPI : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_RRRR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_RRRM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_RRRI : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_RRRF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_RRRP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_RRMR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_RRMM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_RRMI : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_RRMF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_RRMP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_RRIR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_RRIM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_RRIF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_RRIP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_RRFR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_RRFM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_RRFI : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_RRFF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_RRFP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_RRPR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_RRPM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_RRPI : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_RRPF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_RRPP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_RMRR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_RMRM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_RMRI : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_RMRF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_RMRP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_RMMR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_RMMI : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_RMMF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_RMMP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_RMIR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_RMIM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_RMIF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_RMIP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_RMFR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_RMFM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_RMFI : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_RMFF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_RMFP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_RMPR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_RMPM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_RMPI : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_RMPF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_RMPP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_RIRR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_RIRM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_RIRF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_RIRP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_RIMR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_RIMM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_RIMF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_RIMP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_RIFR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_RIFM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_RIFF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_RIFP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_RIPR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_RIPM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_RIPF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_RIPP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_RFRR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_RFRM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_RFRI : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_RFRF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_RFRP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_RFMR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_RFMM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_RFMI : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_RFMF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_RFMP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_RFIR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_RFIM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_RFIF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_RFIP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_RFFR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_RFFM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_RFFI : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_RFPR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_RFPM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_RFPI : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_RPRR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_RPRM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_RPRI : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_RPRF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_RPRP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_RPMR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_RPMM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_RPMI : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_RPMF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_RPMP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_RPIR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_RPIM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_RPIF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_RPIP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_RPFR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_RPFM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_RPFI : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_RPPR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_RPPM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_RPPI : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_MRRR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_MRRM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_MRRI : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_MRRF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_MRRP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_MRMR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_MRMM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_MRMI : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_MRMF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_MRMP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_MRIR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_MRIM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_MRIF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_MRIP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_MRFR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_MRFM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_MRFI : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_MRFF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_MRFP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_MRPR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_MRPM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_MRPI : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_MRPF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_MRPP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_MMRR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_MMRM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_MMRI : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_MMRF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_MMRP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_MMMR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_MMMI : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_MMMF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_MMMP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_MMIR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_MMIM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_MMIF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_MMIP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_MMFR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_MMFM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_MMFI : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_MMFF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_MMFP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_MMPR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_MMPM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_MMPI : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_MMPF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_MMPP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_MIRR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_MIRM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_MIRF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_MIRP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_MIMR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_MIMM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_MIMF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_MIMP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_MIFR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_MIFM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_MIFF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_MIFP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_MIPR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_MIPM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_MIPF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_MIPP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_MFRR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_MFRM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_MFRI : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_MFRF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_MFRP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_MFMR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_MFMM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_MFMI : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_MFMF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_MFMP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_MFIR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_MFIM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_MFIF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_MFIP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_MFFR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_MFFM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_MFFI : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_MFPR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_MFPM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_MFPI : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_MPRR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_MPRM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_MPRI : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_MPRF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_MPRP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_MPMR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_MPMM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_MPMI : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_MPMF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_MPMP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_MPIR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_MPIM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_MPIF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_MPIP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_MPFR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_MPFM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_MPFI : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_MPPR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_MPPM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_MPPI : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_FRRR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_FRRM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_FRRI : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_FRRF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_FRRP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_FRMR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_FRMM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_FRMI : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_FRMF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_FRMP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_FRIR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_FRIM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_FRIF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_FRIP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_FRFR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_FRFM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_FRFI : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_FRFF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_FRFP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_FRPR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_FRPM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_FRPI : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_FRPF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_FRPP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_FMRR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_FMRM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_FMRI : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_FMRF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_FMRP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_FMMR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_FMMI : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_FMMF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_FMMP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_FMIR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_FMIM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_FMIF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_FMIP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_FMFR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_FMFM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_FMFI : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_FMFF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_FMFP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_FMPR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_FMPM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_FMPI : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_FMPF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_FMPP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_FIRR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_FIRM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_FIRF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_FIRP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_FIMR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_FIMM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_FIMF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_FIMP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_FIFR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_FIFM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_FIFF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_FIFP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_FIPR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_FIPM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_FIPF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_FIPP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_FFRR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_FFRM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_FFRI : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_FFRF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_FFRP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_FFMR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_FFMM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_FFMI : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_FFMF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_FFMP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_FFIR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_FFIM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_FFIF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_FFIP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_FFFR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_FFFM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_FFFI : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_FFPR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_FFPM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_FFPI : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_FPRR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_FPRM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_FPRI : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_FPRF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_FPRP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_FPMR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_FPMM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_FPMI : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_FPMF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_FPMP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_FPIR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_FPIM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_FPIF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_FPIP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_FPFR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_FPFM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_FPFI : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_FPPR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_FPPM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMUL_FPPI : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULFWD_RRRX : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULFWD_RRMX : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULFWD_RRIX : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULFWD_RRFX : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULFWD_RRPX : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULFWD_RMRX : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULFWD_RMMX : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULFWD_RMIX : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULFWD_RMFX : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULFWD_RMPX : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULFWD_RIRX : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULFWD_RIMX : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULFWD_RIFX : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULFWD_RIPX : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULFWD_RFRX : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULFWD_RFMX : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULFWD_RFIX : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULFWD_RFFX : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULFWD_RFPX : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULFWD_RPRX : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULFWD_RPMX : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULFWD_RPIX : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULFWD_RPFX : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULFWD_RPPX : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULFWD_MRRX : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULFWD_MRMX : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULFWD_MRIX : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULFWD_MRFX : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULFWD_MRPX : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULFWD_MMRX : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULFWD_MMMX : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULFWD_MMIX : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULFWD_MMFX : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULFWD_MMPX : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULFWD_MIRX : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULFWD_MIMX : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULFWD_MIFX : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULFWD_MIPX : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULFWD_MFRX : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULFWD_MFMX : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULFWD_MFIX : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULFWD_MFFX : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULFWD_MFPX : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULFWD_MPRX : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULFWD_MPMX : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULFWD_MPIX : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULFWD_MPFX : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULFWD_MPPX : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULFWD_FRRX : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULFWD_FRMX : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULFWD_FRIX : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULFWD_FRFX : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULFWD_FRPX : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULFWD_FMRX : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULFWD_FMMX : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULFWD_FMIX : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULFWD_FMFX : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULFWD_FMPX : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULFWD_FIRX : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULFWD_FIMX : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULFWD_FIFX : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULFWD_FIPX : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULFWD_FFRX : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULFWD_FFMX : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULFWD_FFIX : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULFWD_FFFX : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULFWD_FFPX : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULFWD_FPRX : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULFWD_FPMX : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULFWD_FPIX : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULFWD_FPFX : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULFWD_FPPX : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULFWD_RRRX : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULFWD_RRMX : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULFWD_RRIX : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULFWD_RRFX : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULFWD_RRPX : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULFWD_RMRX : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULFWD_RMMX : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULFWD_RMIX : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULFWD_RMFX : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULFWD_RMPX : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULFWD_RIRX : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULFWD_RIMX : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULFWD_RIFX : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULFWD_RIPX : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULFWD_RFRX : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULFWD_RFMX : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULFWD_RFIX : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULFWD_RFFX : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULFWD_RFPX : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULFWD_RPRX : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULFWD_RPMX : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULFWD_RPIX : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULFWD_RPFX : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULFWD_RPPX : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULFWD_MRRX : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULFWD_MRMX : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULFWD_MRIX : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULFWD_MRFX : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULFWD_MRPX : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULFWD_MMRX : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULFWD_MMMX : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULFWD_MMIX : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULFWD_MMFX : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULFWD_MMPX : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULFWD_MIRX : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULFWD_MIMX : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULFWD_MIFX : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULFWD_MIPX : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULFWD_MFRX : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULFWD_MFMX : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULFWD_MFIX : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULFWD_MFFX : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULFWD_MFPX : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULFWD_MPRX : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULFWD_MPMX : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULFWD_MPIX : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULFWD_MPFX : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULFWD_MPPX : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULFWD_FRRX : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULFWD_FRMX : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULFWD_FRIX : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULFWD_FRFX : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULFWD_FRPX : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULFWD_FMRX : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULFWD_FMMX : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULFWD_FMIX : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULFWD_FMFX : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULFWD_FMPX : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULFWD_FIRX : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULFWD_FIMX : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULFWD_FIFX : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULFWD_FIPX : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULFWD_FFRX : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULFWD_FFMX : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULFWD_FFIX : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULFWD_FFFX : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULFWD_FFPX : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULFWD_FPRX : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULFWD_FPMX : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULFWD_FPIX : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULFWD_FPFX : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULFWD_FPPX : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULSRA_RRRR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULSRA_RRRM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULSRA_RRRI : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULSRA_RRRF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULSRA_RRRP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULSRA_RRMR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULSRA_RRMM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULSRA_RRMI : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULSRA_RRMF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULSRA_RRMP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULSRA_RRIR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULSRA_RRIM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULSRA_RRIF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULSRA_RRIP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULSRA_RRFR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULSRA_RRFM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULSRA_RRFI : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULSRA_RRFF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULSRA_RRFP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULSRA_RRPR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULSRA_RRPM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULSRA_RRPI : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULSRA_RRPF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULSRA_RRPP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULSRA_RMRR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULSRA_RMRM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULSRA_RMRI : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULSRA_RMRF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULSRA_RMRP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULSRA_RMMR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULSRA_RMMI : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULSRA_RMMF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULSRA_RMMP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULSRA_RMIR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULSRA_RMIM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULSRA_RMIF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULSRA_RMIP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULSRA_RMFR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULSRA_RMFM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULSRA_RMFI : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULSRA_RMFF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULSRA_RMFP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULSRA_RMPR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULSRA_RMPM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULSRA_RMPI : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULSRA_RMPF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULSRA_RMPP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULSRA_RIRR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULSRA_RIRM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULSRA_RIRF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULSRA_RIRP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULSRA_RIMR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULSRA_RIMM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULSRA_RIMF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULSRA_RIMP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULSRA_RIFR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULSRA_RIFM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULSRA_RIFF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULSRA_RIFP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULSRA_RIPR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULSRA_RIPM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULSRA_RIPF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULSRA_RIPP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULSRA_RFRR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULSRA_RFRM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULSRA_RFRI : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULSRA_RFRF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULSRA_RFRP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULSRA_RFMR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULSRA_RFMM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULSRA_RFMI : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULSRA_RFMF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULSRA_RFMP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULSRA_RFIR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULSRA_RFIM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULSRA_RFIF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULSRA_RFIP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULSRA_RFFR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULSRA_RFFM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULSRA_RFFI : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULSRA_RFPR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULSRA_RFPM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULSRA_RFPI : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULSRA_RPRR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULSRA_RPRM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULSRA_RPRI : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULSRA_RPRF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULSRA_RPRP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULSRA_RPMR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULSRA_RPMM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULSRA_RPMI : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULSRA_RPMF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULSRA_RPMP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULSRA_RPIR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULSRA_RPIM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULSRA_RPIF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULSRA_RPIP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULSRA_RPFR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULSRA_RPFM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULSRA_RPFI : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULSRA_RPPR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULSRA_RPPM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULSRA_RPPI : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULSRA_MRRR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULSRA_MRRM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULSRA_MRRI : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULSRA_MRRF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULSRA_MRRP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULSRA_MRMR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULSRA_MRMM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULSRA_MRMI : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULSRA_MRMF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULSRA_MRMP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULSRA_MRIR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULSRA_MRIM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULSRA_MRIF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULSRA_MRIP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULSRA_MRFR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULSRA_MRFM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULSRA_MRFI : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULSRA_MRFF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULSRA_MRFP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULSRA_MRPR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULSRA_MRPM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULSRA_MRPI : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULSRA_MRPF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULSRA_MRPP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULSRA_MMRR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULSRA_MMRM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULSRA_MMRI : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULSRA_MMRF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULSRA_MMRP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULSRA_MMMR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULSRA_MMMI : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULSRA_MMMF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULSRA_MMMP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULSRA_MMIR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULSRA_MMIF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULSRA_MMIP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULSRA_MMFR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULSRA_MMFM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULSRA_MMFI : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULSRA_MMFF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULSRA_MMFP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULSRA_MMPR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULSRA_MMPM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULSRA_MMPI : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULSRA_MMPF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULSRA_MMPP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULSRA_MIRR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULSRA_MIRM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULSRA_MIRF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULSRA_MIRP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULSRA_MIMR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULSRA_MIMM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULSRA_MIMF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULSRA_MIMP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULSRA_MIFR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULSRA_MIFM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULSRA_MIFF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULSRA_MIFP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULSRA_MIPR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULSRA_MIPM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULSRA_MIPF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULSRA_MIPP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULSRA_MFRR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULSRA_MFRM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULSRA_MFRI : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULSRA_MFRF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULSRA_MFRP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULSRA_MFMR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULSRA_MFMM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULSRA_MFMI : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULSRA_MFMF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULSRA_MFMP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULSRA_MFIR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULSRA_MFIM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULSRA_MFIF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULSRA_MFIP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULSRA_MFFR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULSRA_MFFM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULSRA_MFFI : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULSRA_MFPR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULSRA_MFPM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULSRA_MFPI : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULSRA_MPRR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULSRA_MPRM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULSRA_MPRI : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULSRA_MPRF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULSRA_MPRP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULSRA_MPMR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULSRA_MPMM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULSRA_MPMI : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULSRA_MPMF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULSRA_MPMP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULSRA_MPIR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULSRA_MPIM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULSRA_MPIF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULSRA_MPFR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULSRA_MPFM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULSRA_MPFI : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULSRA_MPPR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULSRA_MPPM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULSRA_MPPI : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULSRA_FRRR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULSRA_FRRM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULSRA_FRRI : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULSRA_FRRF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULSRA_FRRP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULSRA_FRMR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULSRA_FRMM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULSRA_FRMI : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULSRA_FRMF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULSRA_FRMP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULSRA_FRIR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULSRA_FRIM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULSRA_FRIF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULSRA_FRIP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULSRA_FRFR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULSRA_FRFM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULSRA_FRFI : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULSRA_FRFF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULSRA_FRFP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULSRA_FRPR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULSRA_FRPM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULSRA_FRPI : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULSRA_FRPF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULSRA_FRPP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULSRA_FMRR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULSRA_FMRM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULSRA_FMRI : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULSRA_FMRF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULSRA_FMRP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULSRA_FMMR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULSRA_FMMI : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULSRA_FMMF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULSRA_FMMP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULSRA_FMIR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULSRA_FMIF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULSRA_FMIP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULSRA_FMFR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULSRA_FMFM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULSRA_FMFI : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULSRA_FMFF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULSRA_FMFP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULSRA_FMPR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULSRA_FMPM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULSRA_FMPI : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULSRA_FMPF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULSRA_FMPP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULSRA_FIRR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULSRA_FIRM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULSRA_FIRF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULSRA_FIRP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULSRA_FIMR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULSRA_FIMM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULSRA_FIMF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULSRA_FIMP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULSRA_FIFR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULSRA_FIFM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULSRA_FIFF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULSRA_FIFP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULSRA_FIPR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULSRA_FIPM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULSRA_FIPF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULSRA_FIPP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULSRA_FFRR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULSRA_FFRM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULSRA_FFRI : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULSRA_FFRF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULSRA_FFRP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULSRA_FFMR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULSRA_FFMM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULSRA_FFMI : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULSRA_FFMF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULSRA_FFMP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULSRA_FFIR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULSRA_FFIM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULSRA_FFIF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULSRA_FFIP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULSRA_FFFR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULSRA_FFFM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULSRA_FFFI : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULSRA_FFPR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULSRA_FFPM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULSRA_FFPI : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULSRA_FPRR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULSRA_FPRM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULSRA_FPRI : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULSRA_FPRF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULSRA_FPRP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULSRA_FPMR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULSRA_FPMM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULSRA_FPMI : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULSRA_FPMF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULSRA_FPMP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULSRA_FPIR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULSRA_FPIM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULSRA_FPIF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULSRA_FPIP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULSRA_FPFR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULSRA_FPFM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULSRA_FPFI : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULSRA_FPPR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULSRA_FPPM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ADDMULSRA_FPPI : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULSRA_RRRR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULSRA_RRRM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULSRA_RRRI : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULSRA_RRRF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULSRA_RRRP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULSRA_RRMR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULSRA_RRMM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULSRA_RRMI : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULSRA_RRMF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULSRA_RRMP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULSRA_RRIR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULSRA_RRIM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULSRA_RRIF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULSRA_RRIP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULSRA_RRFR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULSRA_RRFM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULSRA_RRFI : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULSRA_RRFF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULSRA_RRFP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULSRA_RRPR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULSRA_RRPM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULSRA_RRPI : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULSRA_RRPF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULSRA_RRPP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULSRA_RMRR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULSRA_RMRM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULSRA_RMRI : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULSRA_RMRF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULSRA_RMRP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULSRA_RMMR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULSRA_RMMI : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULSRA_RMMF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULSRA_RMMP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULSRA_RMIR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULSRA_RMIM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULSRA_RMIF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULSRA_RMIP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULSRA_RMFR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULSRA_RMFM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULSRA_RMFI : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULSRA_RMFF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULSRA_RMFP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULSRA_RMPR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULSRA_RMPM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULSRA_RMPI : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULSRA_RMPF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULSRA_RMPP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULSRA_RIRR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULSRA_RIRM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULSRA_RIRF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULSRA_RIRP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULSRA_RIMR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULSRA_RIMM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULSRA_RIMF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULSRA_RIMP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULSRA_RIFR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULSRA_RIFM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULSRA_RIFF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULSRA_RIFP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULSRA_RIPR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULSRA_RIPM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULSRA_RIPF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULSRA_RIPP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULSRA_RFRR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULSRA_RFRM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULSRA_RFRI : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULSRA_RFRF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULSRA_RFRP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULSRA_RFMR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULSRA_RFMM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULSRA_RFMI : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULSRA_RFMF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULSRA_RFMP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULSRA_RFIR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULSRA_RFIM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULSRA_RFIF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULSRA_RFIP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULSRA_RFFR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULSRA_RFFM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULSRA_RFFI : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULSRA_RFPR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULSRA_RFPM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULSRA_RFPI : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULSRA_RPRR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULSRA_RPRM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULSRA_RPRI : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULSRA_RPRF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULSRA_RPRP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULSRA_RPMR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULSRA_RPMM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULSRA_RPMI : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULSRA_RPMF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULSRA_RPMP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULSRA_RPIR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULSRA_RPIM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULSRA_RPIF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULSRA_RPIP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULSRA_RPFR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULSRA_RPFM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULSRA_RPFI : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULSRA_RPPR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULSRA_RPPM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULSRA_RPPI : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULSRA_MRRR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULSRA_MRRM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULSRA_MRRI : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULSRA_MRRF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULSRA_MRRP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULSRA_MRMR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULSRA_MRMM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULSRA_MRMI : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULSRA_MRMF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULSRA_MRMP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULSRA_MRIR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULSRA_MRIM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULSRA_MRIF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULSRA_MRIP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULSRA_MRFR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULSRA_MRFM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULSRA_MRFI : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULSRA_MRFF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULSRA_MRFP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULSRA_MRPR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULSRA_MRPM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULSRA_MRPI : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULSRA_MRPF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULSRA_MRPP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULSRA_MMRR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULSRA_MMRM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULSRA_MMRI : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULSRA_MMRF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULSRA_MMRP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULSRA_MMMR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULSRA_MMMI : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULSRA_MMMF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULSRA_MMMP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULSRA_MMIR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULSRA_MMIF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULSRA_MMIP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULSRA_MMFR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULSRA_MMFM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULSRA_MMFI : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULSRA_MMFF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULSRA_MMFP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULSRA_MMPR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULSRA_MMPM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULSRA_MMPI : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULSRA_MMPF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULSRA_MMPP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULSRA_MIRR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULSRA_MIRM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULSRA_MIRF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULSRA_MIRP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULSRA_MIMR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULSRA_MIMM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULSRA_MIMF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULSRA_MIMP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULSRA_MIFR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULSRA_MIFM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULSRA_MIFF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULSRA_MIFP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULSRA_MIPR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULSRA_MIPM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULSRA_MIPF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULSRA_MIPP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULSRA_MFRR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULSRA_MFRM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULSRA_MFRI : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULSRA_MFRF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULSRA_MFRP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULSRA_MFMR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULSRA_MFMM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULSRA_MFMI : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULSRA_MFMF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULSRA_MFMP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULSRA_MFIR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULSRA_MFIM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULSRA_MFIP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULSRA_MFFR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULSRA_MFFM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULSRA_MFFI : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULSRA_MFPR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULSRA_MFPM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULSRA_MFPI : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULSRA_MPRR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULSRA_MPRM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULSRA_MPRI : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULSRA_MPRF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULSRA_MPRP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULSRA_MPMR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULSRA_MPMM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULSRA_MPMI : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULSRA_MPMF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULSRA_MPMP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULSRA_MPIR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULSRA_MPIM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULSRA_MPIF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULSRA_MPIP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULSRA_MPFR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULSRA_MPFM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULSRA_MPFI : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULSRA_MPPR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULSRA_MPPM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULSRA_MPPI : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULSRA_FRRR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULSRA_FRRM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULSRA_FRRI : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULSRA_FRRF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULSRA_FRRP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULSRA_FRMR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULSRA_FRMM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULSRA_FRMI : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULSRA_FRMF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULSRA_FRMP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULSRA_FRIR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULSRA_FRIM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULSRA_FRIF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULSRA_FRIP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULSRA_FRFR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULSRA_FRFM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULSRA_FRFI : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULSRA_FRFF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULSRA_FRFP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULSRA_FRPR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULSRA_FRPM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULSRA_FRPI : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULSRA_FRPF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULSRA_FRPP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULSRA_FMRR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULSRA_FMRM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULSRA_FMRI : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULSRA_FMRF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULSRA_FMRP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULSRA_FMMR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULSRA_FMMI : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULSRA_FMMF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULSRA_FMMP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULSRA_FMIR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULSRA_FMIF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULSRA_FMIP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULSRA_FMFR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULSRA_FMFM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULSRA_FMFI : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULSRA_FMFF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULSRA_FMFP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULSRA_FMPR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULSRA_FMPM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULSRA_FMPI : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULSRA_FMPF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULSRA_FMPP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULSRA_FIRR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULSRA_FIRM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULSRA_FIRF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULSRA_FIRP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULSRA_FIMR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULSRA_FIMM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULSRA_FIMF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULSRA_FIMP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULSRA_FIFR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULSRA_FIFM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULSRA_FIFF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULSRA_FIFP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULSRA_FIPR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULSRA_FIPM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULSRA_FIPF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULSRA_FIPP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULSRA_FFRR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULSRA_FFRM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULSRA_FFRI : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULSRA_FFRF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULSRA_FFRP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULSRA_FFMR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULSRA_FFMM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULSRA_FFMI : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULSRA_FFMF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULSRA_FFMP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULSRA_FFIR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULSRA_FFIM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULSRA_FFIF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULSRA_FFIP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULSRA_FFFR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULSRA_FFFM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULSRA_FFFI : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULSRA_FFPR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULSRA_FFPM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULSRA_FFPI : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULSRA_FPRR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULSRA_FPRM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULSRA_FPRI : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULSRA_FPRF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULSRA_FPRP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULSRA_FPMR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULSRA_FPMM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULSRA_FPMI : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULSRA_FPMF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULSRA_FPMP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULSRA_FPIR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULSRA_FPIM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULSRA_FPIF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULSRA_FPIP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULSRA_FPFR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULSRA_FPFM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULSRA_FPFI : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULSRA_FPPR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULSRA_FPPM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SUBMULSRA_FPPI : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ABSDIFF_RXRR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ABSDIFF_RXRM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ABSDIFF_RXRI : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ABSDIFF_RXRF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ABSDIFF_RXRP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ABSDIFF_RXMR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ABSDIFF_RXMM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ABSDIFF_RXMI : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ABSDIFF_RXMF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ABSDIFF_RXMP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ABSDIFF_RXIR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ABSDIFF_RXIM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ABSDIFF_RXIF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ABSDIFF_RXIP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ABSDIFF_RXFR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ABSDIFF_RXFM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ABSDIFF_RXFI : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ABSDIFF_RXFF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ABSDIFF_RXFP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ABSDIFF_RXPR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ABSDIFF_RXPM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ABSDIFF_RXPI : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ABSDIFF_RXPF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ABSDIFF_RXPP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ABSDIFF_MXRR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ABSDIFF_MXRM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ABSDIFF_MXRI : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ABSDIFF_MXRF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ABSDIFF_MXRP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ABSDIFF_MXMR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ABSDIFF_MXMM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ABSDIFF_MXMI : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ABSDIFF_MXMF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ABSDIFF_MXMP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ABSDIFF_MXIR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ABSDIFF_MXIM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ABSDIFF_MXIF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ABSDIFF_MXIP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ABSDIFF_MXFR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ABSDIFF_MXFM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ABSDIFF_MXFI : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ABSDIFF_MXFF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ABSDIFF_MXFP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ABSDIFF_MXPR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ABSDIFF_MXPM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ABSDIFF_MXPI : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ABSDIFF_MXPF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ABSDIFF_MXPP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ABSDIFF_FXRR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ABSDIFF_FXRM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ABSDIFF_FXRI : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ABSDIFF_FXRF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ABSDIFF_FXRP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ABSDIFF_FXMR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ABSDIFF_FXMM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ABSDIFF_FXMI : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ABSDIFF_FXMF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ABSDIFF_FXMP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ABSDIFF_FXIR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ABSDIFF_FXIM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ABSDIFF_FXIF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ABSDIFF_FXIP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ABSDIFF_FXFR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ABSDIFF_FXFM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ABSDIFF_FXFI : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ABSDIFF_FXFF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ABSDIFF_FXFP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ABSDIFF_FXPR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ABSDIFF_FXPM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ABSDIFF_FXPI : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ABSDIFF_FXPF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ABSDIFF_FXPP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ABSDIFFACCUM_RXRR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ABSDIFFACCUM_RXRM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ABSDIFFACCUM_RXRI : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ABSDIFFACCUM_RXRF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ABSDIFFACCUM_RXRP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ABSDIFFACCUM_RXMR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ABSDIFFACCUM_RXMM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ABSDIFFACCUM_RXMI : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ABSDIFFACCUM_RXMF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ABSDIFFACCUM_RXMP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ABSDIFFACCUM_RXIR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ABSDIFFACCUM_RXIM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ABSDIFFACCUM_RXIF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ABSDIFFACCUM_RXIP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ABSDIFFACCUM_RXFR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ABSDIFFACCUM_RXFM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ABSDIFFACCUM_RXFI : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ABSDIFFACCUM_RXFF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ABSDIFFACCUM_RXFP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ABSDIFFACCUM_RXPR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ABSDIFFACCUM_RXPM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ABSDIFFACCUM_RXPI : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ABSDIFFACCUM_RXPF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ABSDIFFACCUM_RXPP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ABSDIFFACCUM_MXRR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ABSDIFFACCUM_MXRM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ABSDIFFACCUM_MXRI : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ABSDIFFACCUM_MXRF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ABSDIFFACCUM_MXRP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ABSDIFFACCUM_MXMR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ABSDIFFACCUM_MXMM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ABSDIFFACCUM_MXMI : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ABSDIFFACCUM_MXMF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ABSDIFFACCUM_MXMP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ABSDIFFACCUM_MXIR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ABSDIFFACCUM_MXIM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ABSDIFFACCUM_MXIF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ABSDIFFACCUM_MXIP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ABSDIFFACCUM_MXFR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ABSDIFFACCUM_MXFM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ABSDIFFACCUM_MXFI : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ABSDIFFACCUM_MXFF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ABSDIFFACCUM_MXFP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ABSDIFFACCUM_MXPR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ABSDIFFACCUM_MXPM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ABSDIFFACCUM_MXPI : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ABSDIFFACCUM_MXPF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ABSDIFFACCUM_MXPP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ABSDIFFACCUM_FXRR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ABSDIFFACCUM_FXRM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ABSDIFFACCUM_FXRI : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ABSDIFFACCUM_FXRF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ABSDIFFACCUM_FXRP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ABSDIFFACCUM_FXMR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ABSDIFFACCUM_FXMM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ABSDIFFACCUM_FXMI : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ABSDIFFACCUM_FXMF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ABSDIFFACCUM_FXMP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ABSDIFFACCUM_FXIR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ABSDIFFACCUM_FXIM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ABSDIFFACCUM_FXIF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ABSDIFFACCUM_FXIP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ABSDIFFACCUM_FXFR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ABSDIFFACCUM_FXFM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ABSDIFFACCUM_FXFI : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ABSDIFFACCUM_FXFF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ABSDIFFACCUM_FXFP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ABSDIFFACCUM_FXPR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ABSDIFFACCUM_FXPM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ABSDIFFACCUM_FXPI : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ABSDIFFACCUM_FXPF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ABSDIFFACCUM_FXPP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ABSDIFFACCUM_XXRR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ABSDIFFACCUM_XXRM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ABSDIFFACCUM_XXRI : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ABSDIFFACCUM_XXRF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ABSDIFFACCUM_XXRP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ABSDIFFACCUM_XXMR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ABSDIFFACCUM_XXMM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ABSDIFFACCUM_XXMI : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ABSDIFFACCUM_XXMF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ABSDIFFACCUM_XXMP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ABSDIFFACCUM_XXIR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ABSDIFFACCUM_XXIM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ABSDIFFACCUM_XXIF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ABSDIFFACCUM_XXIP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ABSDIFFACCUM_XXFR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ABSDIFFACCUM_XXFM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ABSDIFFACCUM_XXFI : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ABSDIFFACCUM_XXFF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ABSDIFFACCUM_XXFP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ABSDIFFACCUM_XXPR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ABSDIFFACCUM_XXPM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ABSDIFFACCUM_XXPI : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ABSDIFFACCUM_XXPF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ABSDIFFACCUM_XXPP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant GET_RXXF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant GET_MXXF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant GET_IXXF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant DECONST_RXXR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant DECONST_RXXM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant DECONST_RXXI : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant DECONST_RXXF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant DECONST_RXXP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant DECONST_MXXR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant DECONST_MXXM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant DECONST_MXXI : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant DECONST_MXXF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant DECONST_MXXP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant DECONST_FXXR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant DECONST_FXXM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant DECONST_FXXI : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant DECONST_FXXF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant DECONST_FXXP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant LDSORT_XXXR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant LDSORT_XXXM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant LDSORT_XXXI : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant LDSORT_XXXF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant LDSORT_XXXP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant UNLDSORT_RXXX : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant UNLDSORT_MXXX : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant UNLDSORT_FXXX : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant CLR_RXXX : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant CLR_IXXX : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant CLR_MXXX : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant CLR_FXXX : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant PUT_FXXR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant PUT_FXXM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant PUT_FXXI : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant PUT_FXXF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant PUT_FXXP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant CMP_XXRR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant CMP_XXRM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant CMP_XXRI : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant CMP_XXRF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant CMP_XXRP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant CMP_XXMR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant CMP_XXMM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant CMP_XXMI : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant CMP_XXMF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant CMP_XXMP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant CMP_XXIR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant CMP_XXIM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant CMP_XXIF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant CMP_XXIP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant CMP_XXFR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant CMP_XXFM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant CMP_XXFI : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant CMP_XXFF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant CMP_XXFP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant CMP_XXPR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant CMP_XXPM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant CMP_XXPI : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant CMP_XXPF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant CMP_XXPP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SETMASKLT_XXRR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SETMASKLT_XXRM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SETMASKLT_XXRI : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SETMASKLT_XXRF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SETMASKLT_XXRP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SETMASKLT_XXMR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SETMASKLT_XXMM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SETMASKLT_XXMI : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SETMASKLT_XXMF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SETMASKLT_XXMP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SETMASKLT_XXIR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SETMASKLT_XXIM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SETMASKLT_XXIF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SETMASKLT_XXIP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SETMASKLT_XXFR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SETMASKLT_XXFM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SETMASKLT_XXFI : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SETMASKLT_XXFF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SETMASKLT_XXFP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SETMASKLT_XXPR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SETMASKLT_XXPM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SETMASKLT_XXPI : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SETMASKLT_XXPF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SETMASKLT_XXPP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SETMASKGT_XXRR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SETMASKGT_XXRM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SETMASKGT_XXRI : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SETMASKGT_XXRF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SETMASKGT_XXRP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SETMASKGT_XXMR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SETMASKGT_XXMM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SETMASKGT_XXMI : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SETMASKGT_XXMF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SETMASKGT_XXMP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SETMASKGT_XXIR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SETMASKGT_XXIM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SETMASKGT_XXIF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SETMASKGT_XXIP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SETMASKGT_XXFR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SETMASKGT_XXFM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SETMASKGT_XXFI : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SETMASKGT_XXFF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SETMASKGT_XXFP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SETMASKGT_XXPR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SETMASKGT_XXPM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SETMASKGT_XXPI : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SETMASKGT_XXPF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SETMASKGT_XXPP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SETMASKEQ_XXRR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SETMASKEQ_XXRM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SETMASKEQ_XXRI : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SETMASKEQ_XXRF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SETMASKEQ_XXRP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SETMASKEQ_XXMR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SETMASKEQ_XXMM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SETMASKEQ_XXMI : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SETMASKEQ_XXMF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SETMASKEQ_XXMP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SETMASKEQ_XXIR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SETMASKEQ_XXIM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SETMASKEQ_XXIF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SETMASKEQ_XXIP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SETMASKEQ_XXFR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SETMASKEQ_XXFM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SETMASKEQ_XXFI : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SETMASKEQ_XXFF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SETMASKEQ_XXFP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SETMASKEQ_XXPR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SETMASKEQ_XXPM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SETMASKEQ_XXPI : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SETMASKEQ_XXPF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SETMASKEQ_XXPP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SETMASKGE_XXRR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SETMASKGE_XXRM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SETMASKGE_XXRI : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SETMASKGE_XXRF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SETMASKGE_XXRP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SETMASKGE_XXMR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SETMASKGE_XXMM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SETMASKGE_XXMI : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SETMASKGE_XXMF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SETMASKGE_XXMP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SETMASKGE_XXIR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SETMASKGE_XXIM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SETMASKGE_XXIF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SETMASKGE_XXIP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SETMASKGE_XXFR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SETMASKGE_XXFM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SETMASKGE_XXFI : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SETMASKGE_XXFF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SETMASKGE_XXFP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SETMASKGE_XXPR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SETMASKGE_XXPM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SETMASKGE_XXPI : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SETMASKGE_XXPF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SETMASKGE_XXPP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SETMASKLE_XXRR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SETMASKLE_XXRM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SETMASKLE_XXRI : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SETMASKLE_XXRF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SETMASKLE_XXRP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SETMASKLE_XXMR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SETMASKLE_XXMM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SETMASKLE_XXMI : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SETMASKLE_XXMF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SETMASKLE_XXMP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SETMASKLE_XXIR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SETMASKLE_XXIM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SETMASKLE_XXIF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SETMASKLE_XXIP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SETMASKLE_XXFR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SETMASKLE_XXFM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SETMASKLE_XXFI : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SETMASKLE_XXFF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SETMASKLE_XXFP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SETMASKLE_XXPR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SETMASKLE_XXPM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SETMASKLE_XXPI : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SETMASKLE_XXPF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SETMASKLE_XXPP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SETMASKNE_XXRR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SETMASKNE_XXRM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SETMASKNE_XXRI : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SETMASKNE_XXRF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SETMASKNE_XXRP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SETMASKNE_XXMR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SETMASKNE_XXMM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SETMASKNE_XXMI : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SETMASKNE_XXMF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SETMASKNE_XXMP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SETMASKNE_XXIR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SETMASKNE_XXIM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SETMASKNE_XXIF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SETMASKNE_XXIP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SETMASKNE_XXFR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SETMASKNE_XXFM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SETMASKNE_XXFI : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SETMASKNE_XXFF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SETMASKNE_XXFP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SETMASKNE_XXPR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SETMASKNE_XXPM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SETMASKNE_XXPI : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SETMASKNE_XXPF : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SETMASKNE_XXPP : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant CMPFWD_XXRX : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant CMPFWD_XXMX : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant CMPFWD_XXIX : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant CMPFWD_XXFX : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant CMPFWD_XXPX : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant PUTFWD_FXXX : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant BARRIERM : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant BARRIERS : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant RPT : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant BEQ : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant BGT : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant BLT : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant BGE : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant BLE : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant BNE : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant INCRXIDXBY1 : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant RESETRXIDX : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant INCTXIDXBY1 : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant RESETTXIDX : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SETSMWB_0 : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant INCSMRB_0 : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant INCSMWB_0 : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SETDMRB_M0 : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SETDMRB_M1 : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SETDMRB_N0 : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SETDMRB_N1 : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SETDMWB_0 : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SETDMWB_1 : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant INCDMRB_M0 : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant INCDMRB_M1 : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant INCDMRB_ALL : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant INCDMRB_N0 : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant INCDMRB_N1 : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant INCDMWB_0 : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant INCDMWB_1 : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant ABSDIFFCLR : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant SORT : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
  constant PUTCA_FXXX : std_logic_vector(3 downto 0) := std_logic_vector(to_unsigned(15, 4));
end;