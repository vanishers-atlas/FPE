library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.std_logic_unsigned.all;

entity testbench is

end entity;

architecture arch of testbench is
	signal 	clock : std_logic := '0';
	signal	kickoff : std_logic := '0';
	signal	running : std_logic;

	signal	PUT_FIFO_0_data  : std_logic_vector(39 downto 0);
	signal	PUT_FIFO_0_write : std_logic;
	signal  PUT_FIFO_0_index : integer := 0;
	type  PUT_FIFO_0_data_array is array (0 to 351) of std_logic_vector(39 downto 0);
	constant PUT_FIFO_0_test_data : PUT_FIFO_0_data_array :=
	(
		-- Test MOV and ACC persistances
		"0000000000000000000000000000000000000000", "0000000000000000000000000000000000000000",
		"0000000000000000000011111111111111111111", "0000000000000000000011111111111111111111",
		"1111111111111111111100000000000000000000", "1111111111111111111100000000000000000000",
		"1111111111111111111111111111111111111111", "1111111111111111111111111111111111111111",

		-- Test LSH 1
		"0010001000100010001000100010001000100010", "0100010001000100010001000100010001000100",
		"1000100010001000100010001000100010001000", "0001000100010001000100010001000100010000",
		"0100010001000100010001000100010001000100", "1000100010001000100010001000100010001000",
		"0001000100010001000100010001000100010000", "0010001000100010001000100010001000100000",
		"1000100010001000100010001000100010001000", "0001000100010001000100010001000100010000",
		"0010001000100010001000100010001000100000", "0100010001000100010001000100010001000000",
		"0001000100010001000100010001000100010000", "0010001000100010001000100010001000100000",
		"0100010001000100010001000100010001000000", "1000100010001000100010001000100010000000",

		-- Test LSH 2
		"0100010001000100010001000100010001000100", "0001000100010001000100010001000100010000",
		"0100010001000100010001000100010001000000", "0001000100010001000100010001000100000000",
		"1000100010001000100010001000100010001000", "0010001000100010001000100010001000100000",
		"1000100010001000100010001000100010000000", "0010001000100010001000100010001000000000",
		"0001000100010001000100010001000100010000", "0100010001000100010001000100010001000000",
		"0001000100010001000100010001000100000000", "0100010001000100010001000100010000000000",
		"0010001000100010001000100010001000100000", "1000100010001000100010001000100010000000",
		"0010001000100010001000100010001000000000", "1000100010001000100010001000100000000000",

		-- Test LSH 3
		"1000100010001000100010001000100010001000", "0100010001000100010001000100010001000000",
		"0010001000100010001000100010001000000000", "0001000100010001000100010001000000000000",
		"0001000100010001000100010001000100010000", "1000100010001000100010001000100010000000",
		"0100010001000100010001000100010000000000", "0010001000100010001000100010000000000000",
		"0010001000100010001000100010001000100000", "0001000100010001000100010001000100000000",
		"1000100010001000100010001000100000000000", "0100010001000100010001000100000000000000",
		"0100010001000100010001000100010001000000", "0010001000100010001000100010001000000000",
		"0001000100010001000100010001000000000000", "1000100010001000100010001000000000000000",

		-- Test LRL 1
		"0010001000100010001000100010001000100010", "0100010001000100010001000100010001000100",
		"1000100010001000100010001000100010001000", "0001000100010001000100010001000100010001",
		"0100010001000100010001000100010001000100", "1000100010001000100010001000100010001000",
		"0001000100010001000100010001000100010001", "0010001000100010001000100010001000100010",
		"1000100010001000100010001000100010001000", "0001000100010001000100010001000100010001",
		"0010001000100010001000100010001000100010", "0100010001000100010001000100010001000100",
		"0001000100010001000100010001000100010001", "0010001000100010001000100010001000100010",
		"0100010001000100010001000100010001000100", "1000100010001000100010001000100010001000",

		-- Test LRL 2
		"0100010001000100010001000100010001000100", "0001000100010001000100010001000100010001",
		"0100010001000100010001000100010001000100", "0001000100010001000100010001000100010001",
		"1000100010001000100010001000100010001000", "0010001000100010001000100010001000100010",
		"1000100010001000100010001000100010001000", "0010001000100010001000100010001000100010",
		"0001000100010001000100010001000100010001", "0100010001000100010001000100010001000100",
		"0001000100010001000100010001000100010001", "0100010001000100010001000100010001000100",
		"0010001000100010001000100010001000100010", "1000100010001000100010001000100010001000",
		"0010001000100010001000100010001000100010", "1000100010001000100010001000100010001000",

		-- Test LRL 3
		"1000100010001000100010001000100010001000", "0100010001000100010001000100010001000100",
		"0010001000100010001000100010001000100010", "0001000100010001000100010001000100010001",
		"0001000100010001000100010001000100010001", "1000100010001000100010001000100010001000",
		"0100010001000100010001000100010001000100", "0010001000100010001000100010001000100010",
		"0010001000100010001000100010001000100010", "0001000100010001000100010001000100010001",
		"1000100010001000100010001000100010001000", "0100010001000100010001000100010001000100",
		"0100010001000100010001000100010001000100", "0010001000100010001000100010001000100010",
		"0001000100010001000100010001000100010001", "1000100010001000100010001000100010001000",

		-- Test RSH 1
		"1100010001000100010001000100010001000100", "1110001000100010001000100010001000100010",
		"1111000100010001000100010001000100010001", "1111100010001000100010001000100010001000",
		"0010001000100010001000100010001000100010", "0001000100010001000100010001000100010001",
		"0000100010001000100010001000100010001000", "0000010001000100010001000100010001000100",
		"0001000100010001000100010001000100010001", "0000100010001000100010001000100010001000",
		"0000010001000100010001000100010001000100", "0000001000100010001000100010001000100010",
		"0000100010001000100010001000100010001000", "0000010001000100010001000100010001000100",
		"0000001000100010001000100010001000100010", "0000000100010001000100010001000100010001",

		-- Test RSH 2
		"1110001000100010001000100010001000100010", "1111100010001000100010001000100010001000",
		"1111111000100010001000100010001000100010", "1111111110001000100010001000100010001000",
		"0001000100010001000100010001000100010001", "0000010001000100010001000100010001000100",
		"0000000100010001000100010001000100010001", "0000000001000100010001000100010001000100",
		"0000100010001000100010001000100010001000", "0000001000100010001000100010001000100010",
		"0000000010001000100010001000100010001000", "0000000000100010001000100010001000100010",
		"0000010001000100010001000100010001000100", "0000000100010001000100010001000100010001",
		"0000000001000100010001000100010001000100", "0000000000010001000100010001000100010001",

		-- Test RSH 3
		"1111000100010001000100010001000100010001", "1111111000100010001000100010001000100010",
		"1111111111000100010001000100010001000100", "1111111111111000100010001000100010001000",
		"0000100010001000100010001000100010001000", "0000000100010001000100010001000100010001",
		"0000000000100010001000100010001000100010", "0000000000000100010001000100010001000100",
		"0000010001000100010001000100010001000100", "0000000010001000100010001000100010001000",
		"0000000000010001000100010001000100010001", "0000000000000010001000100010001000100010",
		"0000001000100010001000100010001000100010", "0000000001000100010001000100010001000100",
		"0000000000001000100010001000100010001000", "0000000000000001000100010001000100010001",

		-- Test RRL 1
		"0100010001000100010001000100010001000100", "0010001000100010001000100010001000100010",
		"0001000100010001000100010001000100010001", "1000100010001000100010001000100010001000",
		"0010001000100010001000100010001000100010", "0001000100010001000100010001000100010001",
		"1000100010001000100010001000100010001000", "0100010001000100010001000100010001000100",
		"0001000100010001000100010001000100010001", "1000100010001000100010001000100010001000",
		"0100010001000100010001000100010001000100", "0010001000100010001000100010001000100010",
		"1000100010001000100010001000100010001000", "0100010001000100010001000100010001000100",
		"0010001000100010001000100010001000100010", "0001000100010001000100010001000100010001",

		-- Test RRL 2
		"0010001000100010001000100010001000100010", "1000100010001000100010001000100010001000",
		"0010001000100010001000100010001000100010", "1000100010001000100010001000100010001000",
		"0001000100010001000100010001000100010001", "0100010001000100010001000100010001000100",
		"0001000100010001000100010001000100010001", "0100010001000100010001000100010001000100",
		"1000100010001000100010001000100010001000", "0010001000100010001000100010001000100010",
		"1000100010001000100010001000100010001000", "0010001000100010001000100010001000100010",
		"0100010001000100010001000100010001000100", "0001000100010001000100010001000100010001",
		"0100010001000100010001000100010001000100", "0001000100010001000100010001000100010001",

		-- Test RRL 3
		"0001000100010001000100010001000100010001", "0010001000100010001000100010001000100010",
		"0100010001000100010001000100010001000100", "1000100010001000100010001000100010001000",
		"1000100010001000100010001000100010001000", "0001000100010001000100010001000100010001",
		"0010001000100010001000100010001000100010", "0100010001000100010001000100010001000100",
		"0100010001000100010001000100010001000100", "1000100010001000100010001000100010001000",
		"0001000100010001000100010001000100010001", "0010001000100010001000100010001000100010",
		"0010001000100010001000100010001000100010", "0100010001000100010001000100010001000100",
		"1000100010001000100010001000100010001000", "0001000100010001000100010001000100010001",

		-- Test NOT
		"1111111111111111111111111111111111111111", "0000000000000000000000000000000000000000",
		"1111111111111111111100000000000000000000", "0000000000000000000011111111111111111111",
		"0000000000000000000011111111111111111111", "1111111111111111111100000000000000000000",
		"0000000000000000000000000000000000000000", "1111111111111111111111111111111111111111",

		-- Test AND
		"0000000000000000000000000000000000000000", "0000000000000000000000000000000000000000", "0000000000000000000000000000000000000000", "1111111111111111111111111111111111111111",
		"0000000000000000000000000000000000000000", "0000000000000000000000000000000000000000", "0000000000000000000000000000000000000000", "1111111111111111111111111111111111111111",
		"0000000000000000000000000000000000000000", "0000000000000000000000000000000000000000", "0000000000000000000000000000000000000000", "1111111111111111111111111111111111111111",
		"0000000000000000000000000000000000000000", "0000000000000000000000000000000000000000", "1111111111111111111111111111111111111111", "1111111111111111111111111111111111111111",

		-- Test NAND
		"1111111111111111111111111111111111111111", "1111111111111111111111111111111111111111", "1111111111111111111111111111111111111111", "0000000000000000000000000000000000000000",
		"1111111111111111111111111111111111111111", "1111111111111111111111111111111111111111", "1111111111111111111111111111111111111111", "0000000000000000000000000000000000000000",
		"1111111111111111111111111111111111111111", "1111111111111111111111111111111111111111", "1111111111111111111111111111111111111111", "0000000000000000000000000000000000000000",
		"1111111111111111111111111111111111111111", "1111111111111111111111111111111111111111", "0000000000000000000000000000000000000000", "0000000000000000000000000000000000000000",

		-- Test OR
		"0000000000000000000000000000000000000000", "1111111111111111111111111111111111111111", "1111111111111111111111111111111111111111", "1111111111111111111111111111111111111111",
		"0000000000000000000000000000000000000000", "1111111111111111111111111111111111111111", "1111111111111111111111111111111111111111", "1111111111111111111111111111111111111111",
		"0000000000000000000000000000000000000000", "1111111111111111111111111111111111111111", "1111111111111111111111111111111111111111", "1111111111111111111111111111111111111111",
		"0000000000000000000000000000000000000000", "0000000000000000000000000000000000000000", "1111111111111111111111111111111111111111", "1111111111111111111111111111111111111111",

		-- Test NOR
		"1111111111111111111111111111111111111111", "0000000000000000000000000000000000000000", "0000000000000000000000000000000000000000", "0000000000000000000000000000000000000000",
		"1111111111111111111111111111111111111111", "0000000000000000000000000000000000000000", "0000000000000000000000000000000000000000", "0000000000000000000000000000000000000000",
		"1111111111111111111111111111111111111111", "0000000000000000000000000000000000000000", "0000000000000000000000000000000000000000", "0000000000000000000000000000000000000000",
		"1111111111111111111111111111111111111111", "1111111111111111111111111111111111111111", "0000000000000000000000000000000000000000", "0000000000000000000000000000000000000000",

		-- Test XOR
		"0000000000000000000000000000000000000000", "1111111111111111111111111111111111111111", "1111111111111111111111111111111111111111", "0000000000000000000000000000000000000000",
		"0000000000000000000000000000000000000000", "1111111111111111111111111111111111111111", "1111111111111111111111111111111111111111", "0000000000000000000000000000000000000000",
		"0000000000000000000000000000000000000000", "1111111111111111111111111111111111111111", "1111111111111111111111111111111111111111", "0000000000000000000000000000000000000000",
		"0000000000000000000000000000000000000000", "0000000000000000000000000000000000000000", "0000000000000000000000000000000000000000", "0000000000000000000000000000000000000000",

		-- Test XNOR
		"1111111111111111111111111111111111111111", "0000000000000000000000000000000000000000", "0000000000000000000000000000000000000000", "1111111111111111111111111111111111111111",
		"1111111111111111111111111111111111111111", "0000000000000000000000000000000000000000", "0000000000000000000000000000000000000000", "1111111111111111111111111111111111111111",
		"1111111111111111111111111111111111111111", "0000000000000000000000000000000000000000", "0000000000000000000000000000000000000000", "1111111111111111111111111111111111111111",
		"1111111111111111111111111111111111111111", "1111111111111111111111111111111111111111", "1111111111111111111111111111111111111111", "1111111111111111111111111111111111111111",

		-- Test ADD
		"0000000000000000000000000000000000000000", "0000000000000000000000000000000000000010",
		"1111111111111111111111111111111111111111", "0000000000000000000000000000000000000000",

		"0000000000000000000000000000000000000000", "0000000000000000000000000000000000000010",
		"1111111111111111111111111111111111111111", "0000000000000000000000000000000000000000",

		"0000000000000000000000000000000000000000", "0000000000000000000000000000000000000010",
		"1111111111111111111111111111111111111111", "0000000000000000000000000000000000000000",

		"0000000000000000000000000000000000000000", "0000000000000000000000000000000000000010",
		"1100110011001100110011001100110011001100", "1111111111111111111111111111111111111110",

		-- Test SUB
		"0000000000000000000000000000000000000010", "0000000000000000000000000000000000000000",
		"1111111111111111111111111111111111111111", "0000000000000000000000000000000000000000",

		"0000000000000000000000000000000000000010", "0000000000000000000000000000000000000000",
		"1111111111111111111111111111111111111111", "0000000000000000000000000000000000000000",

		"0000000000000000000000000000000000000010", "0000000000000000000000000000000000000000",
		"1111111111111111111111111111111111111111", "0000000000000000000000000000000000000000",

		"0000000000000000000000000000000000000000", "0000000000000000000000000000000000000000",
		"0000000000000000000000000000000000000000", "0000000000000000000000000000000000000000",

		-- Test MUL
		"0000000000000000000000000000000000000000", "0000000000000000000000000000000000000000",
		"0000000000000000000000000000000000000001", "0000000000000000000011111110111100000001",

		"0000000000000000000000000000000000000000", "0000000000000000000000000000000000000000",
		"0000000000000000000000000000000000000001", "0000000000000000000011111110111100000001",

		"0000000000000000000000000000000000000000", "0000000000000000000000000000000000000000",
		"0000000000000000000000000000000000000001", "0000000000000000000011111110111100000001",

		"0000000000000000000000000000000000000000", "0000000000000000000000000000000000000001",
		"0000000000000000000000000000000000000100", "0000000000000000000000001111111000000001"

	);

begin
  UUT : entity work.test_FPE_inst(arch)
		port map (
		  PUT_FIFO_0_data  => PUT_FIFO_0_data,
			PUT_FIFO_0_write => PUT_FIFO_0_write,
			clock => clock,
			kickoff => kickoff,
			running => running
		);

  -- Clock generate process
  process
  begin
    loop
      clock <= not clock;
      wait for 50 ns;
    end loop;
  end process;

  -- Signal kickoff after 250 ns
  kickoff <= '1' after 250 ns, '0' after 350 ns;

	-- Check output
	process (clock)
	begin
		if rising_edge(clock) and PUT_FIFO_0_write = '1' then
			-- Check expecting output
			assert(0 <= PUT_FIFO_0_index and PUT_FIFO_0_index < PUT_FIFO_0_test_data'Length)
				report "Unexpected output"
				severity error;

			-- Check the data is correct
			assert(PUT_FIFO_0_data = PUT_FIFO_0_test_data(PUT_FIFO_0_index))
				report "Incorrect " & integer'Image(PUT_FIFO_0_index) & "th output" & lf & ""
				& integer'Image(to_integer(unsigned(PUT_FIFO_0_data))) & " != " & integer'Image(to_integer(unsigned(PUT_FIFO_0_test_data(PUT_FIFO_0_index))))
				severity error;
			assert(PUT_FIFO_0_data /= PUT_FIFO_0_test_data(PUT_FIFO_0_index))
				report "Correct " & integer'Image(PUT_FIFO_0_index) & "th output" & lf & ""
				& integer'Image(to_integer(unsigned(PUT_FIFO_0_data))) & " = " & integer'Image(to_integer(unsigned(PUT_FIFO_0_test_data(PUT_FIFO_0_index))))
				severity note;

			-- Advance to output index
			PUT_FIFO_0_index <= PUT_FIFO_0_index + 1;
		end if;
	end process;

	-- Check end state
	process
	begin
		-- Wait until the end of simulation
		wait for 150 us;

		-- Check all expected output was received
		assert(PUT_FIFO_0_index  = PUT_FIFO_0_test_data'Length)
			report "Not all expected output received"
			severity error;
		assert(PUT_FIFO_0_index /= PUT_FIFO_0_test_data'Length)
			report "all expected output received"
			severity note;
	end process;

end architecture;
